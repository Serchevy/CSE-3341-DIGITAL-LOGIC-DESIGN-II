module MODES
(
	input KEY2, 
	output MODE
);


endmodule 