//module IU 
//(
//	input CLK, RST, 
//	input [3:0] ROW, 
//	output logic [3:0] COL, 
//	output logic [15:0] Input
//);
//	
//	logic [15:0] keyPad;
//	
//	keypad_input INPUT
//	( 
//		.clk(CLK),
//		.reset(RST),
//		.row(ROW),
//		.col(COL),
//		.out(Input)
//	);
//	
//endmodule 